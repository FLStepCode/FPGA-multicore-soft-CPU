`ifndef _noc_parameters_svh_
`define _noc_parameters_svh_

`define PL 33// length of datapack
`define CS 2 // size of single coordinate part
`define RN 9 // number of routers in network

`endif
