`ifndef _queue_parameters_svh_
`define _queue_parameters_svh_

`include "mesh_3x3/inc/noc.svh"

`define EN 4 // number of queue entries
`define EN_B 2 // number of bits required to encode queue entries

`endif
