`define LOAD_REQUESTED  3'b001
`define LOAD_SATISFIED  3'b101
`define STORE_TO_RAM    3'b010