`define TLAST_PRESENT
`define TSTRB_PRESENT