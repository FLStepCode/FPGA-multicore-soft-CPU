// TODO Not actually implemented
module moduleName #(
    parameters
) (
    ports
);
  axis_if_mux;  
endmodule