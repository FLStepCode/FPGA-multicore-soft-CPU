`ifndef _noc_XY_parameters_svh_
`define _noc_XY_parameters_svh_

`define X 3 // number of routers in network on X axis
`define Y 3 // number of routers in network on Y axis

`endif
