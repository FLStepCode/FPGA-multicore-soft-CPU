`ifndef _router_parameters_svh_
`define _router_parameters_svh_

`include "mesh_4x4/inc/noc.svh"

`define REN 5 // number of router entries
`define REN_B 3 // number bits required to eoncode router entries

`endif
