`ifndef _XY_svh_
`define _XY_svh_

`define X 4 // number of routers in network on X axis
`define Y 4 // number of routers in network on Y axis

`endif